module alaw_coder(input_lin, output_alaw);

input [7:0] input_lin;
output [7:0] output_alaw;

endmodule

