module alaw_decoder(input_alaw, output_lin);

input [7:0] input_alaw;
output [7:0] output_lin;

always @(input_alaw) begin
    // TODO: A-law decoder algorithm goes here ;)
end

endmodule

