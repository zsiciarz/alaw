module alaw_coder;

endmodule

